GENERATOR
Time = 0 | rst=0 | d=1 | q=0
DRIVER
Time = 5 | rst=0 | d=1 | q=0
rst = 1
MONITOR
Time = 5 | rst=1 | d=0 | q=0
SCOREBOARD
Time = 5 | rst=1 | d=0 | q=0
-------PASS------
GENERATOR
Time = 5 | rst=0 | d=0 | q=0
MONITOR
Time = 15 | rst=1 | d=1 | q=0
DRIVER
Time = 15 | rst=0 | d=0 | q=0
rst = 1
SCOREBOARD
Time = 15 | rst=1 | d=1 | q=0
-------PASS------
GENERATOR
Time = 15 | rst=0 | d=1 | q=0
MONITOR
Time = 25 | rst=1 | d=0 | q=0
DRIVER
Time = 25 | rst=0 | d=1 | q=0
rst = 1
SCOREBOARD
Time = 25 | rst=1 | d=0 | q=0
-------PASS------
GENERATOR
Time = 25 | rst=0 | d=1 | q=0
MONITOR
Time = 35 | rst=0 | d=1 | q=1
DRIVER
Time = 35 | rst=0 | d=1 | q=0
rst = 0
SCOREBOARD
Time = 35 | rst=0 | d=1 | q=1
-------PASS------
GENERATOR
Time = 35 | rst=0 | d=1 | q=0
MONITOR
Time = 45 | rst=0 | d=1 | q=1
DRIVER
Time = 45 | rst=0 | d=1 | q=0
rst = 0
SCOREBOARD
Time = 45 | rst=0 | d=1 | q=1
-------PASS------

GENERATOR
Time=0  wr=0  d_in=236  addr=11  d_out=0
DRIVER
Time=0  wr=0  d_in=236  addr=11  d_out=0
MONITOR
Time=5  wr=0  d_in=236  addr=11  d_out=0
SCOREBOARD
Time=5  wr=0  d_in=236  addr=11  d_out=0
Read Pass: addr=11 d_out=0
------------------------------------------
GENERATOR
Time=5  wr=0  d_in=184  addr=2  d_out=0
DRIVER
Time=5  wr=0  d_in=184  addr=2  d_out=0
MONITOR
Time=15  wr=0  d_in=184  addr=2  d_out=0
SCOREBOARD
Time=15  wr=0  d_in=184  addr=2  d_out=0
Read Pass: addr=2 d_out=0
------------------------------------------
GENERATOR
Time=15  wr=1  d_in=26  addr=15  d_out=0
DRIVER
Time=15  wr=1  d_in=26  addr=15  d_out=0
MONITOR
Time=25  wr=1  d_in=26  addr=15  d_out=0
SCOREBOARD
Time=25  wr=1  d_in=26  addr=15  d_out=0
Write Pass: addr=15  d_in=26
------------------------------------------
GENERATOR
Time=25  wr=0  d_in=158  addr=9  d_out=0
DRIVER
Time=25  wr=0  d_in=158  addr=9  d_out=0
MONITOR
Time=35  wr=0  d_in=158  addr=9  d_out=0
SCOREBOARD
Time=35  wr=0  d_in=158  addr=9  d_out=0
Read Pass: addr=9 d_out=0
------------------------------------------
GENERATOR
Time=35  wr=1  d_in=167  addr=14  d_out=0
DRIVER
Time=35  wr=1  d_in=167  addr=14  d_out=0
MONITOR
Time=45  wr=1  d_in=167  addr=14  d_out=0
SCOREBOARD
Time=45  wr=1  d_in=167  addr=14  d_out=0
Write Pass: addr=14  d_in=167
------------------------------------------
GENERATOR
Time=45  wr=1  d_in=21  addr=3  d_out=0
DRIVER
Time=45  wr=1  d_in=21  addr=3  d_out=0
MONITOR
Time=55  wr=1  d_in=21  addr=3  d_out=0
SCOREBOARD
Time=55  wr=1  d_in=21  addr=3  d_out=0
Write Pass: addr=3  d_in=21
------------------------------------------
GENERATOR
Time=55  wr=1  d_in=163  addr=3  d_out=0
DRIVER
Time=55  wr=1  d_in=163  addr=3  d_out=0
MONITOR
Time=65  wr=1  d_in=163  addr=3  d_out=0
SCOREBOARD
Time=65  wr=1  d_in=163  addr=3  d_out=0
Write Pass: addr=3  d_in=163
------------------------------------------
GENERATOR
Time=65  wr=1  d_in=53  addr=3  d_out=0
DRIVER
Time=65  wr=1  d_in=53  addr=3  d_out=0
MONITOR
Time=75  wr=1  d_in=53  addr=3  d_out=0
SCOREBOARD
Time=75  wr=1  d_in=53  addr=3  d_out=0
Write Pass: addr=3  d_in=53
------------------------------------------
GENERATOR
Time=75  wr=0  d_in=114  addr=15  d_out=0
DRIVER
Time=75  wr=0  d_in=114  addr=15  d_out=0
MONITOR
Time=85  wr=0  d_in=114  addr=15  d_out=11010
SCOREBOARD
Time=85  wr=0  d_in=114  addr=15  d_out=11010
Read Pass: addr=15 d_out=26
------------------------------------------
GENERATOR
Time=85  wr=0  d_in=230  addr=12  d_out=0
DRIVER
Time=85  wr=0  d_in=230  addr=12  d_out=0
MONITOR
Time=95  wr=0  d_in=230  addr=12  d_out=0
SCOREBOARD
Time=95  wr=0  d_in=230  addr=12  d_out=0
Read Pass: addr=12 d_out=0
------------------------------------------
GENERATOR
Time=95  wr=0  d_in=65  addr=2  d_out=0
DRIVER
Time=95  wr=0  d_in=65  addr=2  d_out=0
MONITOR
Time=105  wr=0  d_in=65  addr=2  d_out=0
SCOREBOARD
Time=105  wr=0  d_in=65  addr=2  d_out=0
Read Pass: addr=2 d_out=0
------------------------------------------
GENERATOR
Time=105  wr=1  d_in=157  addr=10  d_out=0
DRIVER
Time=105  wr=1  d_in=157  addr=10  d_out=0
MONITOR
Time=115  wr=1  d_in=157  addr=10  d_out=0
SCOREBOARD
Time=115  wr=1  d_in=157  addr=10  d_out=0
Write Pass: addr=10  d_in=157
------------------------------------------
GENERATOR
Time=115  wr=1  d_in=18  addr=7  d_out=0
DRIVER
Time=115  wr=1  d_in=18  addr=7  d_out=0
MONITOR
Time=125  wr=1  d_in=18  addr=7  d_out=0
SCOREBOARD
Time=125  wr=1  d_in=18  addr=7  d_out=0
Write Pass: addr=7  d_in=18
------------------------------------------
GENERATOR
Time=125  wr=1  d_in=25  addr=15  d_out=0
DRIVER
Time=125  wr=1  d_in=25  addr=15  d_out=0
MONITOR
Time=135  wr=1  d_in=25  addr=15  d_out=0
SCOREBOARD
Time=135  wr=1  d_in=25  addr=15  d_out=0
Write Pass: addr=15  d_in=25
------------------------------------------
GENERATOR
Time=135  wr=1  d_in=84  addr=5  d_out=0
DRIVER
Time=135  wr=1  d_in=84  addr=5  d_out=0
MONITOR
Time=145  wr=1  d_in=84  addr=5  d_out=0
SCOREBOARD
Time=145  wr=1  d_in=84  addr=5  d_out=0
Write Pass: addr=5  d_in=84
------------------------------------------
GENERATOR
Time=145  wr=1  d_in=66  addr=9  d_out=0
DRIVER
Time=145  wr=1  d_in=66  addr=9  d_out=0
MONITOR
Time=155  wr=1  d_in=66  addr=9  d_out=0
SCOREBOARD
Time=155  wr=1  d_in=66  addr=9  d_out=0
Write Pass: addr=9  d_in=66
------------------------------------------
GENERATOR
Time=155  wr=0  d_in=105  addr=13  d_out=0
DRIVER
Time=155  wr=0  d_in=105  addr=13  d_out=0
MONITOR
Time=165  wr=0  d_in=105  addr=13  d_out=0
SCOREBOARD
Time=165  wr=0  d_in=105  addr=13  d_out=0
Read Pass: addr=13 d_out=0
------------------------------------------
GENERATOR
Time=165  wr=0  d_in=141  addr=0  d_out=0
DRIVER
Time=165  wr=0  d_in=141  addr=0  d_out=0
MONITOR
Time=175  wr=0  d_in=141  addr=0  d_out=0
SCOREBOARD
Time=175  wr=0  d_in=141  addr=0  d_out=0
Read Pass: addr=0 d_out=0
------------------------------------------
GENERATOR
Time=175  wr=1  d_in=17  addr=8  d_out=0
DRIVER
Time=175  wr=1  d_in=17  addr=8  d_out=0
MONITOR
Time=185  wr=1  d_in=17  addr=8  d_out=0
SCOREBOARD
Time=185  wr=1  d_in=17  addr=8  d_out=0
Write Pass: addr=8  d_in=17
------------------------------------------
GENERATOR
Time=185  wr=0  d_in=235  addr=12  d_out=0
DRIVER
Time=185  wr=0  d_in=235  addr=12  d_out=0
MONITOR
Time=195  wr=0  d_in=235  addr=12  d_out=0
SCOREBOARD
Time=195  wr=0  d_in=235  addr=12  d_out=0
Read Pass: addr=12 d_out=0
------------------------------------------

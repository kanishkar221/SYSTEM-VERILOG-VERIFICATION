GENERATOR
Time=0 a=1 b=1 c_in=1 sum=0 c_out=0
DRIVER
Time=1 a=1 b=1 c_in=1 sum=0 c_out=0
MONITOR
Time=2 a=1 b=1 c_in=1 sum=1 c_out=1
SCOREBOARD
Time=2 a=1 b=1 c_in=1 sum=1 c_out=1
=================PASS=================
GENERATOR
Time=3 a=1 b=1 c_in=1 sum=0 c_out=0
DRIVER
Time=4 a=1 b=1 c_in=1 sum=0 c_out=0
MONITOR
Time=5 a=1 b=1 c_in=1 sum=1 c_out=1
SCOREBOARD
Time=5 a=1 b=1 c_in=1 sum=1 c_out=1
=================PASS=================
GENERATOR
Time=6 a=1 b=1 c_in=0 sum=0 c_out=0
DRIVER
Time=7 a=1 b=1 c_in=0 sum=0 c_out=0
MONITOR
Time=8 a=1 b=1 c_in=0 sum=0 c_out=1
SCOREBOARD
Time=8 a=1 b=1 c_in=0 sum=0 c_out=1
=================PASS=================
GENERATOR
Time=9 a=1 b=1 c_in=0 sum=0 c_out=0
DRIVER
Time=10 a=1 b=1 c_in=0 sum=0 c_out=0
MONITOR
Time=11 a=1 b=1 c_in=0 sum=0 c_out=1
SCOREBOARD
Time=11 a=1 b=1 c_in=0 sum=0 c_out=1
=================PASS=================
GENERATOR
Time=12 a=0 b=0 c_in=0 sum=0 c_out=0
DRIVER
Time=13 a=0 b=0 c_in=0 sum=0 c_out=0
MONITOR
Time=14 a=0 b=0 c_in=0 sum=0 c_out=0
SCOREBOARD
Time=14 a=0 b=0 c_in=0 sum=0 c_out=0
=================PASS=================

GENERATOR
Time=0  reset=0  enable=1  count=0
MONITOR
Time=5  reset=0  enable=1  count=1
SOREBOARD
Time=5  reset=0  enable=1  count=1
PASS ----> reset=0  enable=1  Actual count=1  Expected count=1
----------------------------------------------------------------
GENERATOR
Time=10  reset=0  enable=1  count=0
DRIVER
Time=10  reset=0  enable=1  count=0
MONITOR
Time=15  reset=0  enable=1  count=2
SOREBOARD
Time=15  reset=0  enable=1  count=2
PASS ----> reset=0  enable=1  Actual count=2  Expected count=2
----------------------------------------------------------------
GENERATOR
Time=20  reset=0  enable=1  count=0
DRIVER
Time=20  reset=0  enable=1  count=0
MONITOR
Time=25  reset=0  enable=1  count=3
SOREBOARD
Time=25  reset=0  enable=1  count=3
PASS ----> reset=0  enable=1  Actual count=3  Expected count=3
----------------------------------------------------------------
GENERATOR
Time=30  reset=0  enable=1  count=0
DRIVER
Time=30  reset=0  enable=1  count=0
MONITOR
Time=35  reset=0  enable=1  count=4
SOREBOARD
Time=35  reset=0  enable=1  count=4
PASS ----> reset=0  enable=1  Actual count=4  Expected count=4
----------------------------------------------------------------
GENERATOR
Time=40  reset=0  enable=0  count=0
DRIVER
Time=40  reset=0  enable=0  count=0
MONITOR
Time=45  reset=0  enable=0  count=4
SOREBOARD
Time=45  reset=0  enable=0  count=4
PASS ----> reset=0  enable=0  Actual count=4  Expected count=4
----------------------------------------------------------------
GENERATOR
Time=50  reset=0  enable=1  count=0
DRIVER
Time=50  reset=0  enable=1  count=0
MONITOR
Time=55  reset=0  enable=1  count=5
SOREBOARD
Time=55  reset=0  enable=1  count=5
PASS ----> reset=0  enable=1  Actual count=5  Expected count=5
----------------------------------------------------------------
GENERATOR
Time=60  reset=0  enable=0  count=0
DRIVER
Time=60  reset=0  enable=0  count=0
MONITOR
Time=65  reset=0  enable=0  count=5
SOREBOARD
Time=65  reset=0  enable=0  count=5
PASS ----> reset=0  enable=0  Actual count=5  Expected count=5
----------------------------------------------------------------
GENERATOR
Time=70  reset=0  enable=1  count=0
DRIVER
Time=70  reset=0  enable=1  count=0
MONITOR
Time=75  reset=0  enable=1  count=6
SOREBOARD
Time=75  reset=0  enable=1  count=6
PASS ----> reset=0  enable=1  Actual count=6  Expected count=6
----------------------------------------------------------------
GENERATOR
Time=80  reset=0  enable=0  count=0
DRIVER
Time=80  reset=0  enable=0  count=0
MONITOR
Time=85  reset=0  enable=0  count=6
SOREBOARD
Time=85  reset=0  enable=0  count=6
PASS ----> reset=0  enable=0  Actual count=6  Expected count=6
----------------------------------------------------------------
GENERATOR
Time=90  reset=0  enable=1  count=0
DRIVER
Time=90  reset=0  enable=1  count=0
MONITOR
Time=95  reset=0  enable=1  count=7
SOREBOARD
Time=95  reset=0  enable=1  count=7
PASS ----> reset=0  enable=1  Actual count=7  Expected count=7
----------------------------------------------------------------

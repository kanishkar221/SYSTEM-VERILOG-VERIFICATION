GENERATOR
Time=0  rst_n=0  w_en=0  r_en=0  data_in=11101100  data_out=0  full=0  empty=0
MONITOR
Time=5  rst_n=0  w_en=0  r_en=0  data_in=0  data_out=0  full=0  empty=1
SCOREBOARD
Time=5  rst_n=0  w_en=0  r_en=0  data_in=0  data_out=0  full=0  empty=1
RESET : FIFO pointers cleared
----------------------------------------------------------------------------------
GENERATOR
Time=10  rst_n=0  w_en=1  r_en=0  data_in=10111000  data_out=0  full=0  empty=0
DRIVER
Time=10  rst_n=0  w_en=1  r_en=0  data_in=10111000  data_out=0  full=0  empty=0
MONITOR
Time=15  rst_n=1  w_en=1  r_en=0  data_in=10111000  data_out=0  full=0  empty=0
SCOREBOARD
Time=15  rst_n=1  w_en=1  r_en=0  data_in=10111000  data_out=0  full=0  empty=0
WRITE PASS ----> Data written = 184 at location 0
-------------------------------------------------------------------------------------
GENERATOR
Time=20  rst_n=0  w_en=1  r_en=0  data_in=11010  data_out=0  full=0  empty=0
DRIVER
Time=20  rst_n=0  w_en=1  r_en=0  data_in=11010  data_out=0  full=0  empty=0
MONITOR
Time=25  rst_n=1  w_en=1  r_en=0  data_in=11010  data_out=0  full=0  empty=0
SCOREBOARD
Time=25  rst_n=1  w_en=1  r_en=0  data_in=11010  data_out=0  full=0  empty=0
WRITE PASS ----> Data written = 26 at location 1
-------------------------------------------------------------------------------------
GENERATOR
Time=30  rst_n=0  w_en=1  r_en=0  data_in=10011110  data_out=0  full=0  empty=0
DRIVER
Time=30  rst_n=0  w_en=1  r_en=0  data_in=10011110  data_out=0  full=0  empty=0
MONITOR
Time=35  rst_n=1  w_en=1  r_en=0  data_in=10011110  data_out=0  full=0  empty=0
SCOREBOARD
Time=35  rst_n=1  w_en=1  r_en=0  data_in=10011110  data_out=0  full=0  empty=0
WRITE PASS ----> Data written = 158 at location 2
-------------------------------------------------------------------------------------
GENERATOR
Time=40  rst_n=0  w_en=0  r_en=1  data_in=10100111  data_out=0  full=0  empty=0
DRIVER
Time=40  rst_n=0  w_en=0  r_en=1  data_in=10100111  data_out=0  full=0  empty=0
MONITOR
Time=45  rst_n=1  w_en=0  r_en=1  data_in=10100111  data_out=10111000  full=0  empty=0
SCOREBOARD
Time=45  rst_n=1  w_en=0  r_en=1  data_in=10100111  data_out=10111000  full=0  empty=0
READ PASS ----> Actual=184  Expected=184
-------------------------------------------------------------------------------------
GENERATOR
Time=50  rst_n=0  w_en=0  r_en=0  data_in=11100011  data_out=0  full=0  empty=0
DRIVER
Time=50  rst_n=0  w_en=0  r_en=0  data_in=11100011  data_out=0  full=0  empty=0
MONITOR
Time=55  rst_n=1  w_en=0  r_en=0  data_in=11100011  data_out=10111000  full=0  empty=0
SCOREBOARD
Time=55  rst_n=1  w_en=0  r_en=0  data_in=11100011  data_out=10111000  full=0  empty=0
-------------------------------------------------------------------------------------
GENERATOR
Time=60  rst_n=0  w_en=0  r_en=1  data_in=11  data_out=0  full=0  empty=0
DRIVER
Time=60  rst_n=0  w_en=0  r_en=1  data_in=11  data_out=0  full=0  empty=0
MONITOR
Time=65  rst_n=1  w_en=0  r_en=1  data_in=11  data_out=11010  full=0  empty=0
SCOREBOARD
Time=65  rst_n=1  w_en=0  r_en=1  data_in=11  data_out=11010  full=0  empty=0
READ PASS ----> Actual=26  Expected=26
-------------------------------------------------------------------------------------
GENERATOR
Time=70  rst_n=0  w_en=0  r_en=1  data_in=110101  data_out=0  full=0  empty=0
DRIVER
Time=70  rst_n=0  w_en=0  r_en=1  data_in=110101  data_out=0  full=0  empty=0
MONITOR
Time=75  rst_n=1  w_en=0  r_en=1  data_in=110101  data_out=10011110  full=0  empty=1
SCOREBOARD
Time=75  rst_n=1  w_en=0  r_en=1  data_in=110101  data_out=10011110  full=0  empty=1
-------------------------------------------------------------------------------------
GENERATOR
Time=80  rst_n=0  w_en=1  r_en=0  data_in=1110010  data_out=0  full=0  empty=0
DRIVER
Time=80  rst_n=0  w_en=1  r_en=0  data_in=1110010  data_out=0  full=0  empty=0
MONITOR
Time=85  rst_n=1  w_en=1  r_en=0  data_in=1110010  data_out=10011110  full=0  empty=0
SCOREBOARD
Time=85  rst_n=1  w_en=1  r_en=0  data_in=1110010  data_out=10011110  full=0  empty=0
WRITE PASS ----> Data written = 114 at location 3
-------------------------------------------------------------------------------------
GENERATOR
Time=90  rst_n=0  w_en=1  r_en=0  data_in=11100110  data_out=0  full=0  empty=0
DRIVER
Time=90  rst_n=0  w_en=1  r_en=0  data_in=11100110  data_out=0  full=0  empty=0
MONITOR
Time=95  rst_n=1  w_en=1  r_en=0  data_in=11100110  data_out=10011110  full=0  empty=0
SCOREBOARD
Time=95  rst_n=1  w_en=1  r_en=0  data_in=11100110  data_out=10011110  full=0  empty=0
WRITE PASS ----> Data written = 230 at location 4
-------------------------------------------------------------------------------------
